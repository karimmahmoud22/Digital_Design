// Copyright (C) 2023  Intel Corporation. All rights reserved.
// Your use of Intel Corporation's design tools, logic functions 
// and other software and tools, and any partner logic 
// functions, and any output files from any of the foregoing 
// (including device programming or simulation files), and any 
// associated documentation or information are expressly subject 
// to the terms and conditions of the Intel Program License 
// Subscription Agreement, the Intel Quartus Prime License Agreement,
// the Intel FPGA IP License Agreement, or other applicable license
// agreement, including, without limitation, that your use is for
// the sole purpose of programming logic devices manufactured by
// Intel and sold by Intel or its authorized distributors.  Please
// refer to the applicable agreement for further details, at
// https://fpgasoftware.intel.com/eula.

// Generated by Quartus Prime Version 22.1std.2 Build 922 07/20/2023 SC Lite Edition
// Created on Sat Oct 28 11:55:34 2023

// synthesis message_off 10175

`timescale 1ns/1ns

module Assignment (
    reset,clock,W,
    Z);

    input reset;
    input clock;
    input W;
    tri0 reset;
    tri0 W;
    output Z;
    reg Z;
    reg [2:0] fstate;
    reg [2:0] reg_fstate;
    parameter state1=0,state2=1,state3=2;

    always @(posedge clock)
    begin
        if (clock) begin
            fstate <= reg_fstate;
        end
    end

    always @(fstate or reset or W)
    begin
        if (reset) begin
            reg_fstate <= state1;
            Z <= 1'b0;
        end
        else begin
            Z <= 1'b0;
            case (fstate)
                state1: begin
                    if ((W == 1'b1))
                        reg_fstate <= state2;
                    else if ((W == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state1;

                    Z <= 1'b0;
                end
                state2: begin
                    if ((W == 1'b1))
                        reg_fstate <= state3;
                    else if ((W == 1'b0))
                        reg_fstate <= state1;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state2;

                    Z <= 1'b0;
                end
                state3: begin
                    if ((W == 1'b0))
                        reg_fstate <= state1;
                    else if ((W == 1'b1))
                        reg_fstate <= state3;
                    // Inserting 'else' block to prevent latch inference
                    else
                        reg_fstate <= state3;

                    Z <= 1'b1;
                end
                default: begin
                    Z <= 1'bx;
                    $display ("Reach undefined state");
                end
            endcase
        end
    end
endmodule // Assignment
